##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Sat Mar 23 14:31:44 2019
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO rgb2gray
  CLASS BLOCK ;
  SIZE 49.970000 BY 49.980000 ;
  FOREIGN rgb2gray 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.940000 49.910000 29.010000 49.980000 ;
    END
  END clk
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.790000 49.910000 12.860000 49.980000 ;
    END
  END resetn
  PIN r[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 20.390000 49.910000 20.460000 49.980000 ;
    END
  END r[7]
  PIN r[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 19.440000 49.910000 19.510000 49.980000 ;
    END
  END r[6]
  PIN r[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 18.490000 49.910000 18.560000 49.980000 ;
    END
  END r[5]
  PIN r[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 17.540000 49.910000 17.610000 49.980000 ;
    END
  END r[4]
  PIN r[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 16.590000 49.910000 16.660000 49.980000 ;
    END
  END r[3]
  PIN r[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 15.640000 49.910000 15.710000 49.980000 ;
    END
  END r[2]
  PIN r[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 14.690000 49.910000 14.760000 49.980000 ;
    END
  END r[1]
  PIN r[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 13.740000 49.910000 13.810000 49.980000 ;
    END
  END r[0]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.540000 49.910000 36.610000 49.980000 ;
    END
  END b[7]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.590000 49.910000 35.660000 49.980000 ;
    END
  END b[6]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.640000 49.910000 34.710000 49.980000 ;
    END
  END b[5]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.690000 49.910000 33.760000 49.980000 ;
    END
  END b[4]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.740000 49.910000 32.810000 49.980000 ;
    END
  END b[3]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.790000 49.910000 31.860000 49.980000 ;
    END
  END b[2]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.840000 49.910000 30.910000 49.980000 ;
    END
  END b[1]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.890000 49.910000 29.960000 49.980000 ;
    END
  END b[0]
  PIN g[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.990000 49.910000 28.060000 49.980000 ;
    END
  END g[7]
  PIN g[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.040000 49.910000 27.110000 49.980000 ;
    END
  END g[6]
  PIN g[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.090000 49.910000 26.160000 49.980000 ;
    END
  END g[5]
  PIN g[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 25.140000 49.910000 25.210000 49.980000 ;
    END
  END g[4]
  PIN g[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.190000 49.910000 24.260000 49.980000 ;
    END
  END g[3]
  PIN g[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 23.240000 49.910000 23.310000 49.980000 ;
    END
  END g[2]
  PIN g[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.290000 49.910000 22.360000 49.980000 ;
    END
  END g[1]
  PIN g[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 21.340000 49.910000 21.410000 49.980000 ;
    END
  END g[0]
  PIN gray[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 18.490000 0.000000 18.560000 0.070000 ;
    END
  END gray[7]
  PIN gray[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 20.390000 0.000000 20.460000 0.070000 ;
    END
  END gray[6]
  PIN gray[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.290000 0.000000 22.360000 0.070000 ;
    END
  END gray[5]
  PIN gray[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.190000 0.000000 24.260000 0.070000 ;
    END
  END gray[4]
  PIN gray[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.090000 0.000000 26.160000 0.070000 ;
    END
  END gray[3]
  PIN gray[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.990000 0.000000 28.060000 0.070000 ;
    END
  END gray[2]
  PIN gray[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.890000 0.000000 29.960000 0.070000 ;
    END
  END gray[1]
  PIN gray[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.790000 0.000000 31.860000 0.070000 ;
    END
  END gray[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal10 ;
        RECT 46.300000 49.180000 47.100000 49.980000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 46.300000 0.000000 47.100000 0.800000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 2.870000 49.180000 3.670000 49.980000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 2.870000 0.000000 3.670000 0.800000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal10 ;
        RECT 47.900000 49.180000 48.700000 49.980000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 47.900000 0.000000 48.700000 0.800000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 1.270000 49.180000 2.070000 49.980000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 1.270000 0.000000 2.070000 0.800000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 49.970000 49.980000 ;
    LAYER metal2 ;
      RECT 36.680000 49.840000 49.970000 49.980000 ;
      RECT 35.730000 49.840000 36.470000 49.980000 ;
      RECT 34.780000 49.840000 35.520000 49.980000 ;
      RECT 33.830000 49.840000 34.570000 49.980000 ;
      RECT 32.880000 49.840000 33.620000 49.980000 ;
      RECT 31.930000 49.840000 32.670000 49.980000 ;
      RECT 30.980000 49.840000 31.720000 49.980000 ;
      RECT 30.030000 49.840000 30.770000 49.980000 ;
      RECT 29.080000 49.840000 29.820000 49.980000 ;
      RECT 28.130000 49.840000 28.870000 49.980000 ;
      RECT 27.180000 49.840000 27.920000 49.980000 ;
      RECT 26.230000 49.840000 26.970000 49.980000 ;
      RECT 25.280000 49.840000 26.020000 49.980000 ;
      RECT 24.330000 49.840000 25.070000 49.980000 ;
      RECT 23.380000 49.840000 24.120000 49.980000 ;
      RECT 22.430000 49.840000 23.170000 49.980000 ;
      RECT 21.480000 49.840000 22.220000 49.980000 ;
      RECT 20.530000 49.840000 21.270000 49.980000 ;
      RECT 19.580000 49.840000 20.320000 49.980000 ;
      RECT 18.630000 49.840000 19.370000 49.980000 ;
      RECT 17.680000 49.840000 18.420000 49.980000 ;
      RECT 16.730000 49.840000 17.470000 49.980000 ;
      RECT 15.780000 49.840000 16.520000 49.980000 ;
      RECT 14.830000 49.840000 15.570000 49.980000 ;
      RECT 13.880000 49.840000 14.620000 49.980000 ;
      RECT 12.930000 49.840000 13.670000 49.980000 ;
      RECT 0.000000 49.840000 12.720000 49.980000 ;
      RECT 0.000000 0.140000 49.970000 49.840000 ;
      RECT 31.930000 0.000000 49.970000 0.140000 ;
      RECT 30.030000 0.000000 31.720000 0.140000 ;
      RECT 28.130000 0.000000 29.820000 0.140000 ;
      RECT 26.230000 0.000000 27.920000 0.140000 ;
      RECT 24.330000 0.000000 26.020000 0.140000 ;
      RECT 22.430000 0.000000 24.120000 0.140000 ;
      RECT 20.530000 0.000000 22.220000 0.140000 ;
      RECT 18.630000 0.000000 20.320000 0.140000 ;
      RECT 0.000000 0.000000 18.420000 0.140000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 49.970000 49.980000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 49.970000 49.980000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 49.970000 49.980000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 49.970000 49.980000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 49.970000 49.980000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 49.970000 49.980000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 49.970000 49.980000 ;
    LAYER metal10 ;
      RECT 49.500000 48.380000 49.970000 49.980000 ;
      RECT 4.470000 48.380000 45.500000 49.980000 ;
      RECT 0.000000 48.380000 0.470000 49.980000 ;
      RECT 0.000000 1.600000 49.970000 48.380000 ;
      RECT 49.500000 0.000000 49.970000 1.600000 ;
      RECT 4.470000 0.000000 45.500000 1.600000 ;
      RECT 0.000000 0.000000 0.470000 1.600000 ;
  END
END rgb2gray

END LIBRARY
